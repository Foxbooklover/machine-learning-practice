module test;
 initial begin
    $display("Icarus Verilog Test OK!");
    $finish;
  end
endmodule